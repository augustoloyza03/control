library verilog;
use verilog.vl_types.all;
entity control2_vlg_vec_tst is
end control2_vlg_vec_tst;
